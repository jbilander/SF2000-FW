`timescale 1ns / 1ps

module test(
    input a1,
    input a2,
	input a3
);

endmodule
